package common is
    constant common_clk_period : time := 1 ns;
end;
