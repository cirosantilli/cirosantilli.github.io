-- Spaces, tabs and newlines are completely ignored, like C.
-- Semicolons `;` end statements.
-- But indentation and blank lines are nice sometimes.

entity whitespace_tb is end whitespace_tb; architecture behav of whitespace_tb is
begin
process     is
begin
wait; end process;
end behav;
