module display_tb;
    initial
    begin
        $display("hello world");
        $finish;
    end
endmodule
