entity template_tb is
end template_tb;

architecture behav of template_tb is
begin
    process is
    begin
        wait;
    end process;
end behav;
