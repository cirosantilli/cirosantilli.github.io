-- # Comments
--
-- Like this.
--
-- Multiline comments: nope:
-- http://www.thecodingforums.com/threads/multiline-comment.510926/

entity comments_tb is
end entity comments_tb;

architecture behav of comments_tb is
begin
end architecture behav;
