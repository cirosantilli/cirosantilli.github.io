-- Minimal template.

entity min_tb is
end min_tb;

architecture behav of min_tb is
begin
end behav;
